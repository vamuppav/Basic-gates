/home/vamuppav/Documents/ECE637/NOR_pro637/temp/netlist